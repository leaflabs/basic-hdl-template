/*
 * main_zedboard.v
 *
 * Copyright: (C) 2013 LeafLabs, LLC
 * License: MIT License (See LICENSE file)
 * Author: Bryan Newbold <bnewbold@leaflabs.com>
 * Date: November 2013
 *
 */

`timescale 1 ps / 1 ps

module main (
    input wire clock_100mhz,

    // Buttons, LEDs, Switches
    output wire [7:0] leds,
    input wire [7:0] switches,
    input wire button_center,
    input wire button_down,
    input wire button_left,
    input wire button_right,
    input wire button_up,

    // Internal (PS-PL) DDR Interface
    inout wire [15:0] DDR_Addr,
    inout wire [2:0] DDR_BankAddr,
    inout wire DDR_CAS_n,
    inout wire DDR_Clk_n,        // was: DDR_ck_n
    inout wire DDR_Clk_p,        // was: DDR_ck_p
    inout wire DDR_CKE,
    inout wire DDR_CS_n,
    inout wire [3:0] DDR_DM,
    inout wire [31:0] DDR_DQ,
    inout wire [3:0] DDR_DQS_n,
    inout wire [3:0] DDR_DQS_p,
    inout wire DDR_ODT,
    inout wire DDR_RAS_n,
    inout wire DDR_DRSTB,       // was: DDR_reset_n
    inout wire DDR_WEB,         // was: DDR_we_n
    inout wire DDR_VRN,
    inout wire DDR_VRP,

    // Internal (PS-PL) I/O
    inout wire [53:0] MIO,
    inout wire PS_PORB,
    inout wire PS_SRSTB,
    inout wire PS_CLK
    );

    wire axi_aclk;  // This net is the PS's FCLK_CLK0; 100MHz
    wire [0:0] axi_aresetn;
    wire axi_interrupt1;
    wire [31:0] axi_slave1_araddr;
    wire [2:0] axi_slave1_arprot;
    wire [0:0] axi_slave1_arready;
    wire [0:0] axi_slave1_arvalid;
    wire [31:0] axi_slave1_awaddr;
    wire [2:0] axi_slave1_awprot;
    wire [0:0] axi_slave1_awready;
    wire [0:0] axi_slave1_awvalid;
    wire [0:0] axi_slave1_bready;
    wire [1:0] axi_slave1_bresp;
    wire [0:0] axi_slave1_bvalid;
    wire [31:0] axi_slave1_rdata;
    wire [0:0] axi_slave1_rready;
    wire [1:0] axi_slave1_rresp;
    wire [0:0] axi_slave1_rvalid;
    wire [31:0] axi_slave1_wdata;
    wire [0:0] axi_slave1_wready;
    wire [3:0] axi_slave1_wstrb;
    wire [0:0] axi_slave1_wvalid;

    reg throb_led_100mhz = 0;
    reg [25:0] throb_counter_100mhz = 0;
    always @(posedge clock_100mhz) begin
        if (throb_counter_100mhz >= 26'd50_000_000) begin
            throb_counter_100mhz <= 26'd0;
            throb_led_100mhz <= ~throb_led_100mhz;
        end else begin
            throb_counter_100mhz <= throb_counter_100mhz + 26'd1;
        end
    end

    reg throb_led_aclk = 0;
    reg [25:0] throb_counter_aclk = 0;
    always @(posedge axi_aclk) begin
        if (throb_counter_aclk>= 26'd50_000_000) begin
            throb_counter_aclk<= 26'd0;
            throb_led_aclk <= ~throb_led_aclk;
        end else begin
            throb_counter_aclk <= throb_counter_aclk + 26'd1;
        end
    end

    wire [7:0] axi_leds;
    assign leds[0] = axi_leds[0];
    assign leds[1] = axi_leds[1];
    assign leds[2] = axi_leds[2];
    assign leds[3] = axi_leds[3];
    assign leds[4] = button_center;
    assign leds[5] = switches[5];
    assign leds[6] = throb_led_aclk;
    assign leds[7] = throb_led_100mhz;

block_design block_design_i
       (.DDR_addr(DDR_Addr),
        .DDR_ba(DDR_BankAddr),
        .DDR_cas_n(DDR_CAS_n),
        .DDR_ck_n(DDR_Clk_n),
        .DDR_ck_p(DDR_Clk_p),
        .DDR_cke(DDR_CKE),
        .DDR_cs_n(DDR_CS_n),
        .DDR_dm(DDR_DM),
        .DDR_dq(DDR_DQ),
        .DDR_dqs_n(DDR_DQS_n),
        .DDR_dqs_p(DDR_DQS_p),
        .DDR_odt(DDR_ODT),
        .DDR_ras_n(DDR_RAS_n),
        .DDR_reset_n(DDR_DRSTB),
        .DDR_we_n(DDR_WEB),
        .FIXED_IO_ddr_vrn(DDR_VRN),
        .FIXED_IO_ddr_vrp(DDR_VRP),
        .FIXED_IO_mio(MIO),
        .FIXED_IO_ps_clk(PS_CLK),
        .FIXED_IO_ps_porb(PS_PORB),
        .FIXED_IO_ps_srstb(PS_SRSTB),
        .axi_aclk(axi_aclk),
        .axi_aresetn(axi_aresetn),
        .axi_gpio_buttons_tri_i({button_center,
                                 button_down,
                                 button_left,
                                 button_right,
                                 button_up}),
        .axi_gpio_leds_tri_o(axi_leds),
        .axi_interrupt1(axi_interrupt1),
        .axi_slave1_araddr(axi_slave1_araddr),
        .axi_slave1_arprot(axi_slave1_arprot),
        .axi_slave1_arready(axi_slave1_arready),
        .axi_slave1_arvalid(axi_slave1_arvalid),
        .axi_slave1_awaddr(axi_slave1_awaddr),
        .axi_slave1_awprot(axi_slave1_awprot),
        .axi_slave1_awready(axi_slave1_awready),
        .axi_slave1_awvalid(axi_slave1_awvalid),
        .axi_slave1_bready(axi_slave1_bready),
        .axi_slave1_bresp(axi_slave1_bresp),
        .axi_slave1_bvalid(axi_slave1_bvalid),
        .axi_slave1_rdata(axi_slave1_rdata),
        .axi_slave1_rready(axi_slave1_rready),
        .axi_slave1_rresp(axi_slave1_rresp),
        .axi_slave1_rvalid(axi_slave1_rvalid),
        .axi_slave1_wdata(axi_slave1_wdata),
        .axi_slave1_wready(axi_slave1_wready),
        .axi_slave1_wstrb(axi_slave1_wstrb),
        .axi_slave1_wvalid(axi_slave1_wvalid));

axi_lite_slave axi_lite_slave_i (
        .interrupt_request(axi_interrupt1),
        .S_AXI_ACLK(axi_aclk),
        .S_AXI_ARESETN(axi_aresetn),
        .S_AXI_ARADDR(axi_slave1_araddr),
        //.S_AXI_ARPROT(axi_slave1_arprot),
        .S_AXI_ARREADY(axi_slave1_arready),
        .S_AXI_ARVALID(axi_slave1_arvalid),
        .S_AXI_AWADDR(axi_slave1_awaddr),
        //.S_AXI_AWPROT(axi_slave1_awprot),
        .S_AXI_AWREADY(axi_slave1_awready),
        .S_AXI_AWVALID(axi_slave1_awvalid),
        .S_AXI_BREADY(axi_slave1_bready),
        .S_AXI_BRESP(axi_slave1_bresp),
        .S_AXI_BVALID(axi_slave1_bvalid),
        .S_AXI_RDATA(axi_slave1_rdata),
        .S_AXI_RREADY(axi_slave1_rready),
        .S_AXI_RRESP(axi_slave1_rresp),
        .S_AXI_RVALID(axi_slave1_rvalid),
        .S_AXI_WDATA(axi_slave1_wdata),
        .S_AXI_WREADY(axi_slave1_wready),
        .S_AXI_WSTRB(axi_slave1_wstrb),
        .S_AXI_WVALID(axi_slave1_wvalid)
        );
endmodule
